Library IEEE;
Use IEEE.std_logic_1164.all;

Package pBolge is
  Type tBolgeKoord is array(natural range <>) of integer;
End pBolge;
